library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.eig_core_pkg.all;

entity output_loader is

end entity output_loader;

architecture rtl of output_loader is

begin

end architecture rtl;