module tt_um_watchdog 
(
    input  logic clk,
    input  logic rst_n,
    input  logic ena,
    input  logic [7:0] ui_in,       // User Input (7 bits)
    inout wire [7:0] uio,
    output wire [7:0] uio_in,   // Signal, das du aus der Leitung liest
    output wire [7:0] uio_out,  // Signal, das du auf die Leitung schickst
    output wire [7:0] uio_oe    // Steuerung: aktiv für Schreiben (1), Lesen (0)
    output logic [7:0] uo_out      // User Output (8 bits)
);
    logic clk_i;
    logic rst_n_i;
    logic ena_i;

    logic [7:0] ui_in_i;
    logic [7:0] uio_i;
    logic [7:0] uo_out_i;

    // Handshake signals
    logic core_busy_;
    logic res_valid;  // 1-cycle pulse: results ready
    logic ol_busy;
    logic start_ol;
    logic eig_core_start;

    // Data
    logic signed [31:0] alpha, beta;
    logic signed [31:0] invK, K;
    logic [2:0] regime;

    // use bidirectionals as inputs
    // Tri-State Buffer Realisierung
    assign uio = uio_oe ? uio_out : 'z;  // Leitung 'z' wenn lese (uio_oe=0)
    assign uio_in = uio;                  // Lesen immer aufnehmen
    assign clk_i = clk;
    assign ena_i = ena;
    assign rst_n_i = rst_n;
    assign ui_in_i = {1'b0, ui_in};  // Pad ui_in to 8 bits
    assign uio_i = {1'b0, uio_in};    // Pad uio to 8 bits
    assign uo_out = uo_out_i;
        // param_loader Instance
        // Das erzeugst du z.B. so
    initial begin
      uio_out = 8'hA5;  
      uio_oe  = 8'b0;  // Statisch auf 0, Leitung nur lesen
    end
    param_loader u_pl 
    (
        .ena(ena_i),
        .clk(clk_i),
        .rst_n(rst_n),
        .in_pins1(ui_in_i),
        .in_pins2(uio_i),
        .a0(alpha),
        .a1(beta),
        .core_busy(ol_busy && core_busy_),
        .start_calc(eig_core_start)
    );

    // eig_core Instance
    eig_core u_core (
        .ena(ena_i),
        .clk(clk_i),
        .rst_n(rst_n_i),
        .data_rdy(start_ol), 
        .a0(alpha),
        .a1(beta),
        .core_busy(core_busy_),
        .kappa(K),
        .inv_kappa(invK),
        .regime(regime)
    );

    // output_loader Instance
    output_loader u_ol (
        .ena(ena_i),
        .clk(clk_i),
        .rst_n(rst_n_i),
        .start(start_ol),
        .mode(regime),
        .wordA(K),
        .wordB(invK),
        .busy(ol_busy),
        .out_byte(uo_out_i)
    );

always_ff @(posedge clk or negedge rst_n) begin
  if (!rst_n) 
  begin
    //alpha <= 32'b0;
    //beta  <= 32'b0;
    //invK  <= 32'b0;
    //K     <= 32'b0;
    //regime <= 3'b000;
    //uo_out <= 8'b0;
    //core_busy_ <= 1'b0;
    res_valid <= 1'b0;
    //ol_busy <= 1'b0;
    start_ol <= 1'b0;

  end 
  else 
  if (ena) 
  begin 
      eig_core_start <= 1'b1;
      //core_busy_ <= 1'b0;
      //ol_busy <= 1'b0;
  end
  else
  begin
    //uo_out <= 8'b0;
  end
end


endmodule
